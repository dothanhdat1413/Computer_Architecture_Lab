module test_Imm_Gen();
    
endmodule